// FIS types (low byte of the first DWORD)
localparam   FIS_H2DR = 'h27;
localparam   FIS_D2HR = 'h34;
localparam   FIS_DMAA = 'h39;
localparam   FIS_DMAS = 'h41;
localparam   FIS_DATA = 'h46;
localparam   FIS_BIST = 'h58;
localparam   FIS_PIOS = 'h5f;
localparam   FIS_SDB =  'ha1;
