, .INIT_00 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_01 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_02 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_03 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_04 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_05 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_06 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_07 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_08 (256'h2000333040005550555040005550555055505550800080005550800080005550)
, .INIT_09 (256'h19A017401550155019A0155020002AB02490249019A033304000400033303330)
, .INIT_0A (256'h0F1010000BA010001740174012500F10125013B010000E40125013B017401740)
, .INIT_0B (256'h0CD00C300CD00E400AB00CD00BA00AB00B20111015500C300C300C300CD00D80)
, .INIT_0C (256'h0CD00CD013B0174013B00CD01C70333033301C70333040003330400040005550)
, .INIT_0D (256'h0CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD0)
, .INIT_0E (256'h0CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD0)
, .INIT_0F (256'h0CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD00CD0)
