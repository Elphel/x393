// Created with ./create_fold_rom.py
// MCLT 16x16 -> 8x8 fold indices
, .INIT_00 (256'h03A303A203A103A006A806A906AA06AB03B303B203B103B006B806B906BA06BB)
, .INIT_01 (256'h038303820381038006880689068A068B039303920391039006980699069A069B)
, .INIT_02 (256'h001300120011001005180519051A051B000300020001000005080509050A050B)
, .INIT_03 (256'h003300320031003005380539053A053B002300220021002005280529052A052B)
, .INIT_04 (256'h06A406A506A606A70CAF0CAE0CAD0CAC06B406B506B606B70CBF0CBE0CBD0CBC)
, .INIT_05 (256'h06840685068606870C8F0C8E0C8D0C8C06940695069606970C9F0C9E0C9D0C9C)
, .INIT_06 (256'h05140515051605170F1F0F1E0F1D0F1C05040505050605070F0F0F0E0F0D0F0C)
, .INIT_07 (256'h05340535053605370F3F0F3E0F3D0F3C05240525052605270F2F0F2E0F2D0F2C)
, .INIT_08 (256'h0FD30FD20FD10FD00AD80AD90ADA0ADB0FC30FC20FC10FC00AC80AC90ACA0ACB)
, .INIT_09 (256'h0FF30FF20FF10FF00AF80AF90AFA0AFB0FE30FE20FE10FE00AE80AE90AEA0AEB)
, .INIT_0A (256'h036303620361036006680669066A066B037303720371037006780679067A067B)
, .INIT_0B (256'h034303420341034006480649064A064B035303520351035006580659065A065B)
, .INIT_0C (256'h0AD40AD50AD60AD700DF00DE00DD00DC0AC40AC50AC60AC700CF00CE00CD00CC)
, .INIT_0D (256'h0AF40AF50AF60AF700FF00FE00FD00FC0AE40AE50AE60AE700EF00EE00ED00EC)
, .INIT_0E (256'h06640665066606670C6F0C6E0C6D0C6C06740675067606770C7F0C7E0C7D0C7C)
, .INIT_0F (256'h06440645064606470C4F0C4E0C4D0C4C06540655065606570C5F0C5E0C5D0C5C)
