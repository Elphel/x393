, .INIT_00 (256'h000008880FFF0FFF0888044401110111000008880FFF0FFF0888044401110000)
, .INIT_01 (256'h00000222044408880FFF0FFF088808880000044408880FFF0FFF088804440444)
, .INIT_02 (256'h0000000001110222044408880FFF0FFF000001110222044408880FFF0FFF0FFF)
, .INIT_03 (256'h0000000000000000000000000000000000000000000001110222044408880888)
, .INIT_04 (256'h00008888FFFFFFFF888844441111111100008888FFFFFFFF8888444411110000)
, .INIT_05 (256'h0000222244448888FFFFFFFF88888888000044448888FFFFFFFF888844444444)
, .INIT_06 (256'h000000001111222244448888FFFFFFFF00001111222244448888FFFFFFFFFFFF)
, .INIT_07 (256'h0000000000000000000000000000000000000000000011112222444488888888)
