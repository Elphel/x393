/* This is a generated file with the current DDR3 memory timing parameters */

localparam  DLY_LANE0_ODELAY =  80'hd8e8181c1c221c201b20;
localparam  DLY_LANE0_IDELAY =  72'h2078807c88797c7884;
localparam  DLY_LANE1_ODELAY =  80'hd8e31a181b1a1c1c1c1a;
localparam  DLY_LANE1_IDELAY =  72'h247b747b7882787c7c;
localparam          DLY_CMDA = 256'hd4d4d4dadcd3dbd0484848484848484848d4d4ccd4d4dcd9ccd8d4d4d3d3dbd0;
localparam         DLY_PHASE =   8'h32;
// localparam   DFLT_WBUF_DELAY =   4'h8;
