    parameter FPGA_VERSION =          32'h0393003a;