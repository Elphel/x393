// Created with ./create_wnd_mul_rom.py
// MCLT 1d 16 count window with 128:1 super resolution data
, .INIT_00 (256'h0BC80AFF0A36096D08A407DB07110648057F04B603ED0324025B019200C9FFFF)
, .INIT_01 (256'h1857178E16C515FC1533146A13A112D8120F1146107E0FB50EEC0E230D5A0C91)
, .INIT_02 (256'h24E224192351228821BF20F7202E1F651E9D1DD41D0B1C421B7A1AB119E8191F)
, .INIT_03 (256'h3167309F2FD72F0F2E462D7E2CB62BEE2B252A5D299428CC2804273B267325AA)
, .INIT_04 (256'h3DE53D1D3C563B8E3AC639FF3937386F37A736DF3617354F348733BF32F7322F)
, .INIT_05 (256'h4A59499248CB4804473D467645AF44E844204359429241CA4103403C3F743EAC)
, .INIT_06 (256'h56C255FC5536546F53A952E3521C5156508F4FC94F024E3B4D754CAE4BE74B20)
, .INIT_07 (256'h631D6258619360CD60085F425E7D5DB75CF25C2C5B665AA059DA5914584E5788)
, .INIT_08 (256'h6F6A6EA56DE16D1D6C586B946ACF6A0A6946688167BC66F76632656D64A863E3)
, .INIT_09 (256'h7BA57AE17A1E795B789877D47711764D758974C67402733E727A71B670F2702E)
, .INIT_0A (256'h87CC870B8649858784C484028340827D81BB80F880367F737EB07DEE7D2B7C68)
, .INIT_0B (256'h93DF931F925E919E90DD901C8F5B8E9A8DD98D178C568B958AD38A128950888E)
, .INIT_0C (256'h9FDC9F1D9E5D9D9E9CDF9C1F9B609AA099E19921986197A196E19621956094A0)
, .INIT_0D (256'hABBFAB02AA44A986A8C9A80BA74DA68FA5D1A512A454A395A2D7A218A159A09B)
, .INIT_0E (256'hB788B6CCB611B555B498B3DCB320B264B1A7B0EAB02EAF71AEB4ADF7AD3AAC7C)
, .INIT_0F (256'hC335C27BC1C1C107C04CBF92BED8BE1DBD62BCA7BBECBB31BA76B9BBB8FFB844)
, .INIT_10 (256'hCEC4CE0CCD53CC9BCBE3CB2ACA72C9B9C900C847C78EC6D5C61BC562C4A8C3EF)
, .INIT_11 (256'hDA32D97CD8C6D810D75AD6A3D5EDD536D47FD3C8D311D25AD1A2D0EBD033CF7B)
, .INIT_12 (256'hE57FE4CCE418E364E2AFE1FBE146E092DFDDDF28DE73DDBEDD09DC53DB9EDAE8)
, .INIT_13 (256'hF0A9EFF8EF46EE94EDE2ED30EC7EEBCBEB19EA66E9B3E900E84DE79AE6E7E633)
, .INIT_14 (256'hFBAEFAFEFA4FF9A0F8F0F840F790F6E0F630F580F4CFF41FF36EF2BDF20CF15A)
, .INIT_15 (256'h068B05DF0532048503D8032A027D01CF01210074FFC5FF17FE69FDBAFD0CFC5D)
, .INIT_16 (256'h114110970FEC0F420E970DED0D420C960BEB0B400A9409E9093D089107E40738)
, .INIT_17 (256'h1BCC1B241A7D19D5192D188517DD1734168C15E3153A149113E8133E129411EB)
, .INIT_18 (256'h262B258724E2243D239822F2224D21A72101205B1FB51F0E1E681DC11D1A1C73)
, .INIT_19 (256'h305D2FBC2F1A2E772DD52D332C902BED2B4A2AA72A03296028BC2818277426D0)
, .INIT_1A (256'h3A6039C23923388337E4374536A53605356534C53424338332E3324231A030FF)
, .INIT_1B (256'h4433439742FB425F41C34127408A3FED3F503EB33E153D783CDA3C3C3B9D3AFF)
, .INIT_1C (256'h4DD44D3B4CA24C094B704AD74A3D49A4490A487047D5473B46A04605456A44CF)
, .INIT_1D (256'h574156AC5616558054EA545453BE5327529151FA516350CB50344F9C4F044E6C)
, .INIT_1E (256'h60795FE75F555EC35E305D9D5D0A5C775BE45B505ABC5A28599458FF586B57D6)
, .INIT_1F (256'h697B68EC685E67CF674066B0662165916501647163E0635062BF622E619C610B)
, .INIT_20 (256'h724571BA712F70A370186F8C6F006E746DE76D5A6CCD6C406BB36B256A976A09)
, .INIT_21 (256'h7AD67A4F79C7793F78B7782F77A6771E7695760C758274F9746F73E5735A72D0)
, .INIT_22 (256'h832D82A9822581A1811D809880137F8E7F097E837DFD7D777CF17C6B7BE47B5D)
, .INIT_23 (256'h8B488AC88A4889C7894788C6884587C3874286C0863E85BC853984B6843383B0)
, .INIT_24 (256'h932692A9922D91B1913490B7903A8FBC8F3E8EC08E428DC48D458CC68C478BC7)
, .INIT_25 (256'h9AC59A4D99D5995C98E3986A97F1977796FD96839609958E95139498941D93A1)
, .INIT_26 (256'hA226A1B2A13DA0C9A0549FDE9F699EF39E7E9E079D919D1A9CA39C2C9BB59B3D)
, .INIT_27 (256'hA946A8D6A865A7F5A784A713A6A1A630A5BEA54CA4D9A467A3F4A381A30DA29A)
, .INIT_28 (256'hB024AFB8AF4CAEDFAE73AE06AD98AD2BACBDAC4FABE1AB72AB04AA94AA25A9B6)
, .INIT_29 (256'hB6C0B658B5F0B588B51FB4B6B44DB3E4B37AB311B2A6B23CB1D1B166B0FBB090)
, .INIT_2A (256'hBD18BCB4BC51BBEDBB88BB24BABFBA5AB9F4B98FB929B8C3B85CB7F6B78FB727)
, .INIT_2B (256'hC32BC2CCC26DC20DC1ADC14DC0ECC08BC02ABFC9BF67BF05BEA3BE41BDDEBD7B)
, .INIT_2C (256'hC8F9C89EC843C7E8C78CC730C6D4C678C61BC5BEC561C503C4A5C447C3E9C38A)
, .INIT_2D (256'hCE81CE2ACDD4CD7DCD25CCCECC76CC1ECBC6CB6DCB14CABBCA62CA08C9AEC954)
, .INIT_2E (256'hD3C1D36FD31DD2CAD277D224D1D1D17ED12AD0D6D081D02CCFD7CF82CF2DCED7)
, .INIT_2F (256'hD8B9D86BD81ED7D0D782D733D6E4D695D646D5F6D5A6D556D506D4B5D464D412)
, .INIT_30 (256'hDD68DD1FDCD6DC8DDC43DBF9DBAFDB64DB19DACEDA83DA37D9EBD99FD953D906)
, .INIT_31 (256'hE1CDE189E145E100E0BBE075E030DFEADFA4DF5DDF17DECFDE88DE40DDF9DDB0)
, .INIT_32 (256'hE5E8E5A9E569E529E4E9E4A8E467E426E3E4E3A2E360E31EE2DBE298E255E211)
, .INIT_33 (256'hE9B9E97EE943E907E8CCE890E853E817E7DAE79DE75FE722E6E3E6A5E667E628)
, .INIT_34 (256'hED3DED07ECD1EC9AEC63EC2CEBF4EBBDEB84EB4CEB13EADAEAA1EA67EA2DE9F3)
, .INIT_35 (256'hF076F045F013EFE1EFAFEF7CEF4AEF17EEE3EEAFEE7CEE47EE13EDDEEDA9ED73)
, .INIT_36 (256'hF362F336F309F2DCF2AEF281F253F224F1F6F1C7F197F168F138F108F0D8F0A7)
, .INIT_37 (256'hF601F5D9F5B1F589F561F538F50FF4E5F4BBF491F467F43CF411F3E6F3BAF38E)
, .INIT_38 (256'hF853F830F80DF7E9F7C6F7A2F77DF759F734F70EF6E9F6C3F69DF676F650F629)
, .INIT_39 (256'hFA57FA39FA1AF9FCF9DDF9BEF99EF97FF95EF93EF91DF8FCF8DBF8B9F898F875)
, .INIT_3A (256'hFC0DFBF3FBDAFBC0FBA6FB8CFB72FB57FB3BFB20FB04FAE8FACBFAAFFA92FA74)
, .INIT_3B (256'hFD74FD60FD4BFD37FD21FD0CFCF6FCE0FCCAFCB3FC9DFC85FC6EFC56FC3EFC25)
, .INIT_3C (256'hFE8DFE7EFE6EFE5EFE4EFE3EFE2DFE1CFE0AFDF9FDE7FDD4FDC2FDAFFD9BFD88)
, .INIT_3D (256'hFF57FF4DFF42FF37FF2CFF20FF15FF08FEFCFEEFFEE2FED5FEC7FEB9FEAAFE9C)
, .INIT_3E (256'hFFD2FFCDFFC7FFC1FFBBFFB4FFADFFA6FF9FFF97FF8FFF86FF7DFF74FF6BFF61)
, .INIT_3F (256'hFFFFFFFEFFFEFFFDFFFBFFF9FFF7FFF5FFF3FFF0FFECFFE9FFE5FFE1FFDCFFD8)
, .INITP_00 (256'h0000000000000000000000000000000000000000000000000000000000000001)
, .INITP_02 (256'h5555555555555555555550000000000000000000000000000000000000000000)
, .INITP_03 (256'h5555555555555555555555555555555555555555555555555555555555555555)
, .INITP_04 (256'h5555555555555555555555555555555555555555555555555555555555555555)
, .INITP_05 (256'h5555555555555555555555555555555555555555555555555555555555555555)
, .INITP_06 (256'h5555555555555555555555555555555555555555555555555555555555555555)
, .INITP_07 (256'h5555555555555555555555555555555555555555555555555555555555555555)
