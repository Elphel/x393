, .INIT_00 (256'hF1EFE1CED1ADC18CB16BA14A9129810870E760C650A540843063204210210000)
, .INIT_01 (256'hE3DEF3FFC39CD3BDA35AB37B8318933962D672F7429452B52252327302101231)
, .INIT_02 (256'hD58DC5ACF5CFE5EE95098528B54BA56A548544A474C764E61401042034432462)
, .INIT_03 (256'hC7BCD79DE7FEF7DF87389719A77AB75B46B4569566F676D70630161126723653)
, .INIT_04 (256'hB92BA90A99698948F9AFE98ED9EDC9CC382328021861084078A7688658E548C4)
, .INIT_05 (256'hAB1ABB3B8B589B79EB9EFBBFCBDCDBFD2A123A330A501A716A967AB74AD45AF5)
, .INIT_06 (256'h9D498D68BD0BAD2ADDCDCDECFD8FEDAE1C410C603C032C225CC54CE47C876CA6)
, .INIT_07 (256'h8F789F59AF3ABF1BCFFCDFDDEFBEFF9F0E701E512E323E134EF45ED56EB67E97)
, .INIT_08 (256'h606770464025500420E330C200A11080E16FF14EC12DD10CA1EBB1CA81A99188)
, .INIT_09 (256'h725662775214423532D222F3129002B1F35EE37FD31CC33DB3DAA3FB939883B9)
, .INIT_0A (256'h4405542464477466048114A024C334E2C50DD52CE54FF56E858995A8A5CBB5EA)
, .INIT_0B (256'h563446157676665716B0069136F226D3D73CC71DF77EE75F97B88799B7FAA7DB)
, .INIT_0C (256'h28A3388208E118C06827780648655844A9ABB98A89E999C8E92FF90EC96DD94C)
, .INIT_0D (256'h3A922AB31AD00AF17A166A375A544A75BB9AABBB9BD88BF9FB1EEB3FDB5CCB7D)
, .INIT_0E (256'h0CC11CE02C833CA24C455C646C077C268DC99DE8AD8BBDAACD4DDD6CED0FFD2E)
, .INIT_0F (256'h1EF00ED13EB22E935E744E557E366E179FF88FD9BFBAAF9BDF7CCF5DFF3EEF1F)
