/home/andrey/git/x393/includes/x393_cur_params_target_00.vh