, .INITP_00 (INITP_00)
, .INITP_01 (INITP_01)
, .INITP_02 (INITP_02)
, .INITP_03 (INITP_03)
, .INITP_04 (INITP_04)
, .INITP_05 (INITP_05)
, .INITP_06 (INITP_06)
, .INITP_07 (INITP_07)
, .INITP_08 (INITP_08)
, .INITP_09 (INITP_09)
, .INITP_0A (INITP_0A)
, .INITP_0B (INITP_0B)
, .INITP_0C (INITP_0C)
, .INITP_0D (INITP_0D)
, .INITP_0E (INITP_0E)
, .INITP_0F (INITP_0F)
, .INIT_00  (INIT_00)
, .INIT_01  (INIT_01)
, .INIT_02  (INIT_02)
, .INIT_03  (INIT_03)
, .INIT_04  (INIT_04)
, .INIT_05  (INIT_05)
, .INIT_06  (INIT_06)
, .INIT_07  (INIT_07)
, .INIT_08  (INIT_08)
, .INIT_09  (INIT_09)
, .INIT_0A  (INIT_0A)
, .INIT_0B  (INIT_0B)
, .INIT_0C  (INIT_0C)
, .INIT_0D  (INIT_0D)
, .INIT_0E  (INIT_0E)
, .INIT_0F  (INIT_0F)
, .INIT_10  (INIT_10)
, .INIT_11  (INIT_11)
, .INIT_12  (INIT_12)
, .INIT_13  (INIT_13)
, .INIT_14  (INIT_14)
, .INIT_15  (INIT_15)
, .INIT_16  (INIT_16)
, .INIT_17  (INIT_17)
, .INIT_18  (INIT_18)
, .INIT_19  (INIT_19)
, .INIT_1A  (INIT_1A)
, .INIT_1B  (INIT_1B)
, .INIT_1C  (INIT_1C)
, .INIT_1D  (INIT_1D)
, .INIT_1E  (INIT_1E)
, .INIT_1F  (INIT_1F)
, .INIT_20  (INIT_20)
, .INIT_21  (INIT_21)
, .INIT_22  (INIT_22)
, .INIT_23  (INIT_23)
, .INIT_24  (INIT_24)
, .INIT_25  (INIT_25)
, .INIT_26  (INIT_26)
, .INIT_27  (INIT_27)
, .INIT_28  (INIT_28)
, .INIT_29  (INIT_29)
, .INIT_2A  (INIT_2A)
, .INIT_2B  (INIT_2B)
, .INIT_2C  (INIT_2C)
, .INIT_2D  (INIT_2D)
, .INIT_2E  (INIT_2E)
, .INIT_2F  (INIT_2F)
, .INIT_30  (INIT_30)
, .INIT_31  (INIT_31)
, .INIT_32  (INIT_32)
, .INIT_33  (INIT_33)
, .INIT_34  (INIT_34)
, .INIT_35  (INIT_35)
, .INIT_36  (INIT_36)
, .INIT_37  (INIT_37)
, .INIT_38  (INIT_38)
, .INIT_39  (INIT_39)
, .INIT_3A  (INIT_3A)
, .INIT_3B  (INIT_3B)
, .INIT_3C  (INIT_3C)
, .INIT_3D  (INIT_3D)
, .INIT_3E  (INIT_3E)
, .INIT_3F  (INIT_3F)
, .INIT_40  (INIT_40)
, .INIT_41  (INIT_41)
, .INIT_42  (INIT_42)
, .INIT_43  (INIT_43)
, .INIT_44  (INIT_44)
, .INIT_45  (INIT_45)
, .INIT_46  (INIT_46)
, .INIT_47  (INIT_47)
, .INIT_48  (INIT_48)
, .INIT_49  (INIT_49)
, .INIT_4A  (INIT_4A)
, .INIT_4B  (INIT_4B)
, .INIT_4C  (INIT_4C)
, .INIT_4D  (INIT_4D)
, .INIT_4E  (INIT_4E)
, .INIT_4F  (INIT_4F)
, .INIT_50  (INIT_50)
, .INIT_51  (INIT_51)
, .INIT_52  (INIT_52)
, .INIT_53  (INIT_53)
, .INIT_54  (INIT_54)
, .INIT_55  (INIT_55)
, .INIT_56  (INIT_56)
, .INIT_57  (INIT_57)
, .INIT_58  (INIT_58)
, .INIT_59  (INIT_59)
, .INIT_5A  (INIT_5A)
, .INIT_5B  (INIT_5B)
, .INIT_5C  (INIT_5C)
, .INIT_5D  (INIT_5D)
, .INIT_5E  (INIT_5E)
, .INIT_5F  (INIT_5F)
, .INIT_60  (INIT_60)
, .INIT_61  (INIT_61)
, .INIT_62  (INIT_62)
, .INIT_63  (INIT_63)
, .INIT_64  (INIT_64)
, .INIT_65  (INIT_65)
, .INIT_66  (INIT_66)
, .INIT_67  (INIT_67)
, .INIT_68  (INIT_68)
, .INIT_69  (INIT_69)
, .INIT_6A  (INIT_6A)
, .INIT_6B  (INIT_6B)
, .INIT_6C  (INIT_6C)
, .INIT_6D  (INIT_6D)
, .INIT_6E  (INIT_6E)
, .INIT_6F  (INIT_6F)
, .INIT_70  (INIT_70)
, .INIT_71  (INIT_71)
, .INIT_72  (INIT_72)
, .INIT_73  (INIT_73)
, .INIT_74  (INIT_74)
, .INIT_75  (INIT_75)
, .INIT_76  (INIT_76)
, .INIT_77  (INIT_77)
, .INIT_78  (INIT_78)
, .INIT_79  (INIT_79)
, .INIT_7A  (INIT_7A)
, .INIT_7B  (INIT_7B)
, .INIT_7C  (INIT_7C)
, .INIT_7D  (INIT_7D)
, .INIT_7E  (INIT_7E)
, .INIT_7F  (INIT_7F)
