// Created with ./create_wnd_sres4_rom.py
// MCLT 16x16  window with 4:1 super resolution data
, .INIT_00 (256'h238721BE1FE01DEE1BEA19D517AF157C133A10ED0E960C3509CD075F04ED0277)
, .INIT_01 (256'h323F322F320131B4314830BD30152F4F2E6C2D6C2C502B1929C7285B26D7253B)
, .INIT_02 (256'h46F943673FAC3BCA37C3339A2F502AEA266921D01D23186313950EBA09D704ED)
, .INIT_03 (256'h645F644063E363486271615C600C5E815CBB5ABC588556175374509E4D964A5E)
, .INIT_04 (256'h6A3E64E75F525981537A4D3F46D4403E3980329E2B9E24821D50160C0EBA075F)
, .INIT_05 (256'h96409612958794A0935D91C08FC88D788AD087D3848380E07CEE78AF74256F54)
, .INIT_06 (256'h8D4386297EBC77016EFD66B45E2C556A4C73434D39FE308A26F91D50139509CD)
, .INIT_07 (256'hC7C6C788C6CFC59CC3EFC1C9BF2BBC18B891B497B02FAB5AA61BA0759A6D9405)
, .INIT_08 (256'hAFF0A7179DD894378A3B7FEA754A6A615F3753D2483A3C75308A248218630C35)
, .INIT_09 (256'hF8D0F883F79DF61EF408F15BEE19EA44E5DFE0ECDB6ED569CEE1C7D9C055B85B)
, .INIT_0A (256'hD230C79FBC93B112A52598D18C1F7F1771C16424564A483A39FE2B9E1D230E96)
, .INIT_0B (256'h294028E427D22608238A20581C7317E012A00CB60627FEF6F728EEC1E5C7DC3F)
, .INIT_0C (256'hF3EFE7ACDAD9CD80BFA8B15AA29F937F84047438642453D2434D329E21D010ED)
, .INIT_0D (256'h58F9588F5750553D52584EA34A1F44CF3EB737DA303D27E51ED615160AABFF9C)
, .INIT_0E (256'h15170729F899E96FD9B6C976B8B9A78B95F6840471C15F374C7339802669133A)
, .INIT_0F (256'h87DE876585FB83A080567C1F76FE70F66A0A623E5998501D45D33AC02EEB225B)
, .INIT_10 (256'h3595260515BF04CEF33DE115CE62BB31A78B937F7F176A61556A403E2AEA157C)
, .INIT_11 (256'hB5D1B54AB3B5B113AD67A8B2A2F69C39947D8BC8821E77876C085FA8526F4466)
, .INIT_12 (256'h5554442B323A1F8D0C2EF829E38CCE62B8B9A29F8C1F754A5E2C46D42F5017AF)
, .INIT_13 (256'hE2B5E221E062DD7CD96FD43ECDECC67EBDF7B45DA9B69E08915B83B7752365AA)
, .INIT_14 (256'h744061894DF8399924790EA5F829E115C976B15A98D17FEA66B44D3F339A19D5)
, .INIT_15 (256'h0E700DCE0BE708BE0453FEAAF7C5EFAAE65EDBE5D047C38BB5B8A6D796F18611)
, .INIT_16 (256'h92467E0D68E852E53C1124790C2EF33DD9B6BFA8A5258A3B6EFD537A37C31BEA)
, .INIT_17 (256'h38E73837362A32BF2DF827DA206817A50D990248F5BAE7F7D906C8F2B7C4A587)
, .INIT_18 (256'hAF5599A682FA6B5F52E539991F8D04CEE96FCD80B1129437770159813BCA1DEE)
, .INIT_19 (256'h61FE61425F0E5B6456464FB747BA3E563390276E19F70B36FB31E9F4D788C3FA)
, .INIT_1A (256'hCB59B4419C1D82FA68E84DF8323A15BFF899DAD9BC939DD87EBC5F523FAC1FE0)
, .INIT_1B (256'h899E88D5867D82967D2276266DA563A4582B4B3F3CE92D321C2309C7F629E155)
, .INIT_1C (256'hE642CDD0B44199A67E0D6189442B26050729E7ACC79FA717862964E7436721BE)
, .INIT_1D (256'hAFACAED8AC5DA83BA2769B119210877A7B546DA65E794DD63BC828581394FD88)
, .INIT_1E (256'hFFFFE642CB59AF5592467440555435951517F3EFD230AFF08D436A3E46F92387)
, .INIT_1F (256'hD413D334D097CC3DC629BE60B4E5A9C09CF58E8E7E946D0F5A0C45952FB81881)
, .INIT_20 (256'h1881FD88E155C3FAA587861165AA4466225BFF9CDC3FB85B94056F544A5E253B)
, .INIT_21 (256'hF6BBF5D1F314EE85E827DFFED60FCA61BCFAADE29D248AC976DD616B4A82322F)
, .INIT_22 (256'h2FB81394F629D788B7C496F17523526F2EEB0AABE5C7C0559A6D74254D9626D7)
, .INIT_23 (256'h178F169B13C00EFE085AFFD6F57AE94ADB4ECB90BA18A6F292287BC963E24A82)
, .INIT_24 (256'h4595285809C7E9F4C8F2A6D783B75FA83AC01516EEC1C7D9A07578AF509E285B)
, .INIT_25 (256'h367B357E32852D9426AD1DD513110667F7E0E784D55DC177ABDE94A07BC9616B)
, .INIT_26 (256'h5A0C3BC81C23FB31D906B5B8915B6C0845D31ED6F728CEE1A61B7CEE537429C7)
, .INIT_27 (256'h536C52654F524A35431039E82EC221A7129C01ADEEE3DA4AC3EEABDE922876DD)
, .INIT_28 (256'h6D0F4DD62D320B36E7F7C38B9E087787501D27E5FEF6D569AB5A80E056172B19)
, .INIT_29 (256'h6E506D416A1564CE5D6F53FD487E3AF82B7419FC069AF15ADA4AC177A6F28AC9)
, .INIT_2A (256'h7E945E793CE919F7F5BAD047A9B6821E5998303D0627DB6EB02F848358852C50)
, .INIT_2B (256'h871585FF82BC7D4F75BB6C056033524B425730611C73069AEEE3D55DBA189D24)
, .INIT_2C (256'h8E8E6DA64B3F276E0248DBE5B45D8BC8623E37DA0CB6E0ECB49787D35ABC2D6C)
, .INIT_2D (256'h9DAE9C91993993AA8BE581F175D26792573844CE306119FC01ADE784CB90ADE2)
, .INIT_2E (256'h9CF57B54582B33900D99E65EBDF7947D6A0A3EB712A0E5DFB8918AD05CBB2E6C)
, .INIT_2F (256'hB20DB0E9AD7EA7CF9FDF95B289507ABF6A09573842572B74129CF7E0DB4EBCFA)
, .INIT_30 (256'hA9C0877A63A43E5617A5EFAAC67E9C3970F644CF17E0EA44BC188D785E812F4F)
, .INIT_31 (256'hC423C2FABF7FB9B4B19DA73E9A9F8BC77ABF6792524B3AF821A70667E94ACA61)
, .INIT_32 (256'hB4E592106DA547BA2068F7C5CDECA2F676FE4A1F1C73EE19BF2B8FC8600C3015)
, .INIT_33 (256'hD3E7D2B9CF2FC94CC113B689A9B59A9F895075D26033487E2EC21311F57AD60F)
, .INIT_34 (256'hBE609B1176264FB727DAFEAAD43EA8B27C1F4EA32058F15BC1C991C0615C30BD)
, .INIT_35 (256'hE14FE01DDC86D68FCE39C38AB689A73E95B281F16C0553FD39E81DD5FFD6DFFE)
, .INIT_36 (256'hC629A2767D2256462DF80453D96FAD6780565258238AF408C3EF935D62713148)
, .INIT_37 (256'hEC52EB1CE77CE173D906CE39C113B19D9FDF8BE575BB5D6F431026AD085AE827)
, .INIT_38 (256'hCC3DA83B82965B6432BF08BEDD7CB11383A0553D2608F61EC59C94A0634831B4)
, .INIT_39 (256'hF4EAF3B1F009E9F3E173D68FC94CB9B4A7CF93AA7D4F64CE4A352D940EFEEE85)
, .INIT_3A (256'hD097AC5D867D5F0E362A0BE7E062B3B585FB575027D2F79DC6CF958763E33201)
, .INIT_3B (256'hFB11F9D6F628F009E77CDC86CF2FBF7FAD7E993982BC6A154F52328513C0F314)
, .INIT_3C (256'hD334AED888D5614238370DCEE221B54A8765588F28E4F883C78896126440322F)
, .INIT_3D (256'hFEC3FD88F9D6F3B1EB1CE01DD2B9C2FAB0E99C9185FF6D415265357E169BF5D1)
, .INIT_3E (256'hD413AFAC899E61FE38E70E70E2B5B5D187DE58F92940F8D0C7C69640645F323F)
, .INIT_3F (256'hFFFFFEC3FB11F4EAEC52E14FD3E7C423B20D9DAE87156E50536C367B178FF6BB)
, .INITP_01 (256'h5555555550000000555555540000000055555400000000000000000000000000)
, .INITP_02 (256'hAAAAA55555540000AA9555555550000055555555554000005555555555000000)
, .INITP_03 (256'hAAAAAAAA55554000AAAAAAA955554000AAAAAAA555550000AAAAAA5555550000)
, .INITP_04 (256'hFFFFFAAAA9555000FFFFAAAAA9555000FFEAAAAAA5555000AAAAAAAA95554000)
, .INITP_05 (256'hFFFFFFEAAA955400FFFFFFEAAA955400FFFFFFAAAA555400FFFFFEAAAA555000)
, .INITP_06 (256'hFFFFFFFEAAA55400FFFFFFFAAA955400FFFFFFFAAA955400FFFFFFFAAA955400)
, .INITP_07 (256'hFFFFFFFEAAA55400FFFFFFFEAAA55400FFFFFFFEAAA55400FFFFFFFEAAA55400)
