// Created with ./create_wnd_mul_rom.py
// MCLT 1d 16 count window with 128:1 super resolution data
, .INIT_00 (256'h1921178F15FD146B12D911470FB50E230C910AFF096D07DB064804B603240192)
, .INIT_01 (256'h323F30AD2F1B2D8A2BF82A6628D4274325B1241F228D20FB1F691DD71C451AB3)
, .INIT_02 (256'h4B5449C3483246A14510437F41ED405C3ECB3D393BA83A17388536F4356233D0)
, .INIT_03 (256'h645F62CE613E5FAE5E1D5C8D5AFC596C57DB564A54BA5329519850074E764CE5)
, .INIT_04 (256'h7D597BCA7A3B78AB771C758D73FD726E70DE6F4E6DBF6C2F6A9F690F677F65EF)
, .INIT_05 (256'h964094B39325919790098E7A8CEC8B5E89CF884186B285248395820680777EE8)
, .INIT_06 (256'hAF10AD84ABF8AA6BA8DFA752A5C5A439A2ACA11E9F919E049C779AE9995C97CE)
, .INIT_07 (256'hC7C6C63BC4B1C326C19BC010BE85BCFABB6FB9E3B858B6CCB540B3B5B229B09D)
, .INIT_08 (256'hE05CDED3DD4BDBC2DA39D8B0D727D59ED415D28BD102CF78CDEECC64CADAC950)
, .INIT_09 (256'hF8D0F749F5C3F43DF2B6F12FEFA8EE21EC9AEB13E98CE804E67CE4F4E36CE1E4)
, .INIT_0A (256'h111D0F990E150C910B0D09890805068004FB037601F1006CFEE7FD61FBDBFA56)
, .INIT_0B (256'h294027BF263E24BD233B21BA20381EB61D341BB21A2F18AD172A15A7142412A0)
, .INIT_0C (256'h41353FB83E393CBB3B3D39BE383F36C0354133C1324230C22F422DC22C412AC1)
, .INIT_0D (256'h58F9577F56045489530D519250164E9A4D1E4BA14A2548A8472B45AE443142B3)
, .INIT_0E (256'h70886F116D996C216AA9693167B9664064C8634E61D5605C5EE25D685BEE5A74)
, .INIT_0F (256'h87DE866A84F68382820E80997F247DAF7C3A7AC5794F77D9766374EC737671FF)
, .INIT_10 (256'h9EF79D879C179AA7993797C6965594E493729201908F8F1C8DAA8C378AC48951)
, .INIT_11 (256'hB5D1B465B2F9B18DB020AEB4AD47ABDAAA6CA8FEA790A622A4B4A345A1D6A067)
, .INIT_12 (256'hCC66CAFFC998C830C6C8C55FC3F6C28DC124BFBBBE51BCE7BB7DBA12B8A7B73C)
, .INIT_13 (256'hE2B5E153DFEFDE8CDD28DBC5DA60D8FCD797D632D4CDD367D201D09BCF34CDCE)
, .INIT_14 (256'hF8BAF75CF5FDF49FF340F1E1F081EF21EDC1EC61EB00E99FE83EE6DCE57AE418)
, .INIT_15 (256'h0E700D170BBE0A64090A07B0065504FA039F024300E8FF8BFE2FFCD2FB75FA18)
, .INIT_16 (256'h23D62282212E1FD91E841D2F1BDA1A84192E17D71680152913D2127A11220FC9)
, .INIT_17 (256'h38E73798364934FA33AB325B310B2FBA2E692D182BC62A74292227D0267D2529)
, .INIT_18 (256'h4DA04C574B0E49C4487A473045E5449A434F420340B73F6A3E1E3CD03B833A35)
, .INIT_19 (256'h61FE60BB5F785E345CF05BAB5A66592157DB5695554E540752C0517950314EE9)
, .INIT_1A (256'h75FF74C17384724671086FC96E8A6D4A6C0A6ACA698A6849670765C664846341)
, .INIT_1B (256'h899E8867872F85F784BF8387824E81147FDB7EA07D667C2B7AF079B47878773B)
, .INIT_1C (256'h9CD99BA89A779945981496E195AF947B9348921490E08FAB8E768D418C0B8AD4)
, .INIT_1D (256'hAFACAE82AD58AC2DAB01A9D6A8A9A77DA650A522A3F4A2C6A197A0689F399E09)
, .INIT_1E (256'hC216C0F3BFCFBEABBD86BC61BB3BBA15B8EFB7C8B6A1B579B451B328B200B0D6)
, .INIT_1F (256'hD413D2F7D1DAD0BCCF9ECE80CD61CC42CB22CA02C8E2C7C1C6A0C57EC45CC339)
, .INIT_20 (256'hE5A0E48BE375E25EE148E030DF19DE00DCE8DBCFDAB5D99BD881D766D64BD52F)
, .INIT_21 (256'hF6BBF5ADF49EF38FF27FF16FF05FEF4EEE3CED2AEC18EB05E9F2E8DEE7CAE6B5)
, .INIT_22 (256'h0761065A0553044B0343023A01310027FF1DFE12FD07FBFCFAF0F9E3F8D6F7C9)
, .INIT_23 (256'h178F169015901490138F128E118C108A0F870E840D810C7C0B780A73096D0867)
, .INIT_24 (256'h2743264C2554245B23622268216E20741F791E7D1D811C851B881A8A198D188E)
, .INIT_25 (256'h367B358B349B33AA32B931C730D52FE22EEF2DFB2D072C122B1D2A282931283B)
, .INIT_26 (256'h4534444C4364427B419240A83FBE3ED33DE83CFC3C103B233A3539483859376B)
, .INIT_27 (256'h536C528C51AC50CB4FEA4F094E264D444C604B7D4A9849B448CE47E84702461B)
, .INIT_28 (256'h612060495F715E995DC05CE65C0C5B325A57597B589F57C356E55608552A544B)
, .INIT_29 (256'h6E506D816CB16BE16B106A3F696E689B67C966F66622654E647963A462CE61F7)
, .INIT_2A (256'h7AF77A31796A78A277DA77117648757F74B473EA731E7253718670B96FEC6F1E)
, .INIT_2B (256'h87158658859984DA841B835B829A81D9811880557F937ED07E0C7D477C837BBD)
, .INIT_2C (256'h92A891F3913E90888FD18F1A8E628DA98CF18C378B7D8AC28A07894C889087D3)
, .INIT_2D (256'h9DAE9D029C559BA89AFA9A4C999D98ED983D978D96DB962A957794C49411935D)
, .INIT_2E (256'hA826A782A6DFA63AA595A4F0A44AA3A3A2FCA254A1ACA103A05A9FB09F059E5A)
, .INIT_2F (256'hB20DB172B0D8B03CAFA0AF04AE67ADC9AD2BAC8DABEDAB4DAAADAA0CA96AA8C8)
, .INIT_30 (256'hBB62BAD1BA3FB9ADB91AB887B7F3B75EB6C9B634B59EB507B470B3D8B33FB2A6)
, .INIT_31 (256'hC423C39BC313C28AC201C177C0ECC061BFD5BF48BEBBBE2EBDA0BD11BC82BBF2)
, .INIT_32 (256'hCC50CBD2CB53CAD3CA53C9D2C951C8CFC84CC7C9C746C6C1C63CC5B7C531C4AA)
, .INIT_33 (256'hD3E7D372D2FDD286D210D198D120D0A8D02FCFB5CF3ACEC0CE44CDC8CD4BCCCE)
, .INIT_34 (256'hDAE7DA7CDA0FD9A3D935D8C7D859D7EAD77AD70AD699D627D5B5D543D4CFD45C)
, .INIT_35 (256'hE14FE0EDE08AE027DFC3DF5FDEFADE94DE2EDDC7DD60DCF8DC8FDC26DBBCDB52)
, .INIT_36 (256'hE71DE6C5E66CE612E5B8E55DE502E4A6E449E3ECE38EE330E2D1E271E211E1B0)
, .INIT_37 (256'hEC52EC03EBB4EB64EB13EAC2EA70EA1EE9CBE977E923E8CEE879E823E7CCE775)
, .INIT_38 (256'hF0ECF0A7F061F01BEFD4EF8CEF44EEFCEEB2EE68EE1EEDD3ED87ED3BECEEECA0)
, .INIT_39 (256'hF4EAF4AEF472F436F3F9F3BBF37DF33EF2FEF2BEF27DF23CF1FAF1B7F174F130)
, .INIT_3A (256'hF84CF81AF7E8F7B5F782F74EF719F6E4F6AEF678F641F609F5D1F598F55EF524)
, .INIT_3B (256'hFB11FAE9FAC1FA98FA6EFA44FA19F9EEF9C2F995F968F93AF90CF8DCF8ADF87C)
, .INIT_3C (256'hFD39FD1BFCFCFCDDFCBDFC9DFC7CFC5BFC38FC16FBF2FBCEFBA9FB84FB5EFB38)
, .INIT_3D (256'hFEC3FEAFFE9BFE85FE6FFE59FE42FE2AFE12FDF9FDDFFDC5FDAAFD8FFD73FD56)
, .INIT_3E (256'hFFB0FFA6FF9BFF90FF84FF77FF6AFF5CFF4DFF3EFF2FFF1EFF0DFEFCFEE9FED7)
, .INIT_3F (256'hFFFFFFFFFFFEFFFCFFFAFFF7FFF4FFF0FFEBFFE6FFE0FFDAFFD3FFCBFFC3FFBA)
, .INITP_01 (256'h5555555555555555555555555555555555555555555555000000000000000000)
, .INITP_02 (256'hAAAAAAAAAAAAAAAAAAAAA9555555555555555555555555555555555555555555)
, .INITP_03 (256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA)
, .INITP_04 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAA)
, .INITP_05 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INITP_06 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INITP_07 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
