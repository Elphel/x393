, .INIT_00 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_01 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_02 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_03 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_04 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_05 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_06 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_07 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_08 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_09 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_0A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_0B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_0C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_0D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_0E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_0F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_10 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_11 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_12 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_13 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_14 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_15 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_16 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_17 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_18 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_19 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_1A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_1B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_1C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_1D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_1E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_1F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_20 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_21 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_22 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_23 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_24 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_25 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_26 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_27 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_28 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_29 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_2A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_2B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_2C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_2D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_2E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_2F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_30 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_31 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_32 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_33 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_34 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_35 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_36 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_37 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_38 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_39 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_3A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_3B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_3C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_3D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_3E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_3F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_40 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_41 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_42 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_43 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_44 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_45 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_46 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_47 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_48 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_49 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_4A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_4B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_4C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_4D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_4E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_4F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_50 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_51 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_52 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_53 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_54 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_55 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_56 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_57 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_58 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_59 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_5A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_5B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_5C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_5D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_5E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_5F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_60 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_61 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_62 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_63 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_64 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_65 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_66 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_67 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_68 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_69 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_6A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_6B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_6C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_6D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_6E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_6F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
, .INIT_70 (256'h103C103810341030102C102810241020101C101810141010100C100810041000)
, .INIT_71 (256'h107C107810741070106C106810641060105C105810541050104C104810441040)
, .INIT_72 (256'h10BC10B810B410B010AC10A810A410A0109C109810941090108C108810841080)
, .INIT_73 (256'h10FC10F810F410F010EC10E810E410E010DC10D810D410D010CC10C810C410C0)
, .INIT_74 (256'h113C113811341130112C112811241120111C111811141110110C110811041100)
, .INIT_75 (256'h117C117811741170116C116811641160115C115811541150114C114811441140)
, .INIT_76 (256'h11BC11B811B411B011AC11A811A411A0119C119811941190118C118811841180)
, .INIT_77 (256'h11FC11F811F411F011EC11E811E411E011DC11D811D411D011CC11C811C411C0)
, .INIT_78 (256'h123C123812341230122C122812241220121C121812141210120C120812041200)
, .INIT_79 (256'h127C127812741270126C126812641260125C125812541250124C124812441240)
, .INIT_7A (256'h12BC12B812B412B012AC12A812A412A0129C129812941290128C128812841280)
, .INIT_7B (256'h12FC12F812F412F012EC12E812E412E012DC12D812D412D012CC12C812C412C0)
, .INIT_7C (256'h133C133813341330132C132813241320131C131813141310130C130813041300)
, .INIT_7D (256'h137C137813741370136C136813641360135C135813541350134C134813441340)
, .INIT_7E (256'h13BC13B813B413B013AC13A813A413A0139C139813941390138C138813841380)
, .INIT_7F (256'h0FFC13F813F413F013EC13E813E413E013DC13D813D413D013CC13C813C413C0)
