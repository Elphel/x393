// Created with ./create_rotator_rom.py
// MCLT rotator cos/sin values
, .INIT_00 (256'hFFDCFFE5FFECFFF3FFF7FFFBFFFEFFFF0000000000000000000000000000FFFF)
, .INIT_01 (256'hFEC7FF15FF57FF8FFFBBFFDCFFF3FFFEFF74FF97FFB4FFCDFFE1FFF0FFF9FFFE)
, .INIT_02 (256'hFC9DFD74FE2DFEC7FF42FF9FFFDCFFFBFDD4FE5EFED5FF37FF86FFC1FFE9FFFD)
, .INIT_03 (256'hF95EFB04FC6EFD9BFE8DFF42FFBBFFF7FB20FC56FD60FE3EFEEFFF74FFCDFFF9)
, .INIT_04 (256'hF50FF7C6FA1AFC0DFD9BFEC7FF8FFFF3F759F97FFB57FCE0FE1CFF08FFA6FFF5)
, .INIT_05 (256'hEFAFF3BAF734FA1AFC6EFE2DFF57FFECF281F5D9F8B9FB20FD0CFE7EFF74FFF0)
, .INIT_06 (256'hE943EEE3F3BAF7C6FB04FD74FF15FFE5EC9AF168F589F8FCFBC0FDD4FF37FFE9)
, .INIT_07 (256'hE1CDE943EFAFF50FF95EFC9DFEC7FFDCE5A9EC2CF1C7F676FA39FD0CFEEFFFE1)
, .INIT_08 (256'hD953E2DBEB13F1F6F77DFBA6FE6EFFD2DDB0E628ED73F38EF875FC25FE9CFFD8)
, .INIT_09 (256'hCFD7DBAFE5E8EE7CF561FA92FE0AFFC7D4B5DF5DE890F045F676FB20FE3EFFCD)
, .INIT_0A (256'hC561D3C1E030EAA1F309F95EFD9BFFBBCABBD7D0E31EEC9AF43CF9FCFDD4FFC1)
, .INIT_0B (256'hB9F4CB14D9EBE667F076F80DFD21FFADBFC9CF82DD1FE890F1C7F8B9FD60FFB4)
, .INIT_0C (256'hAD98C1ADD31DE1CDEDA9F69DFC9DFF9FB3E4C678D695E426EF17F759FCE0FFA6)
, .INIT_0D (256'hA054B78FCBC6DCD6EAA1F50FFC0DFF8FA713BCB4CF82DF5DEC2CF5D9FC56FF97)
, .INIT_0E (256'h922DACBDC3E9D782E75FF362FB72FF7D995CB23CC7E8DA37E907F43CFBC0FF86)
, .INIT_0F (256'h832DA13DBB88D1D1E3E4F197FACBFF6B8AC8A713BFC9D4B5E5A9F281FB20FF74)
, .INIT_10 (256'h735A9513B2A6CBC6E030EFAFFA1AFF577B5D9B3DB727CED7E211F0A7FA74FF61)
, .INIT_11 (256'h62BF8845A946C561DC43EDA9F95EFF426B258EC0AE06C89EDE40EEAFF9BEFF4D)
, .INIT_12 (256'h51637AD69F69BEA3D81EEB84F898FF2C5A2881A1A467C20DDA37EC9AF8FCFF37)
, .INIT_13 (256'h3F506CCD9513B78FD3C1E943F7C6FF15487073E59A4DBB24D5F6EA67F830FF20)
, .INIT_14 (256'h2C905E308A48B024CF2DE6E3F6E9FEFC360565918FBCB3E4D17EE817F759FF08)
, .INIT_15 (256'h192D4F047F09A865CA62E467F601FEE222F256AC84B6AC4FCCCEE5A9F676FEEF)
, .INIT_16 (256'h05323F50735AA054C561E1CDF50FFEC70F42473B793FA467C7E8E31EF589FED5)
, .INIT_17 (256'hF0A92F1A674097F1C02ADF17F411FEAAFAFE37456D5A9C2CC2CCE075F491FEB9)
, .INIT_18 (256'hDB9E1E685ABC8F3EBABFDC43F309FE8DE63326D0610B93A1BD7BDDB0F38EFE9C)
, .INIT_19 (256'hC61B0D424DD4863EB51FD953F1F6FE6ED0EB15E354548AC8B7F6DACEF281FE7E)
, .INIT_1A (256'hB02EFBAE408A7CF1AF4CD646F0D8FE4EBB310485473B81A1B23CD7D0F168FE5E)
, .INIT_1B (256'h99E1E9B332E3735AA946D31DEFAFFE2DA512F2BD39C2782FAC4FD4B5F045FE3E)
, .INIT_1C (256'h8340D75A24E2697BA30DCFD7EE7CFE0A8E9AE0922BED6E74A630D17EEF17FE1C)
, .INIT_1D (256'h6C58C4A8168C5F559CA3CC76ED3DFDE777D4CE0C1DC164719FDECE2AEDDEFDF9)
, .INIT_1E (256'h5536B1A707E454EA9609C8F9EBF4FDC260CDBB310F425A28995CCABBEC9AFDD4)
, .INIT_1F (256'h3DE59E5DF8F04A3D8F3EC561EAA1FD9B4992A80B00744F9C92A9C730EB4CFDAF)
, .INIT_20 (256'h0BC80A3608A40711057F03ED025B00C9FD88E9F3C38A8BC744CFF15A94A0322F)
, .INIT_21 (256'h23511E9D19E81533107E0BC80711025B178E146A11460E230AFF07DB04B60192)
, .INIT_22 (256'h3AC632F72B2523511B7A13A10BC803ED2F0F28CC22881C4215FC0FB5096D0324)
, .INIT_23 (256'h521C473D3C56316726731B7A107E057F46763D1D33BF2A5D20F7178E0E2304B6)
, .INIT_24 (256'h69465B664D753F7431672351153307115DB7515644E8386F2BEE1F6512D80648)
, .INIT_25 (256'h80366F6A5E7D4D753C562B2519E808A474C6656D55FC467636DF273B178E07DB)
, .INIT_26 (256'h96E183406F6A5B66473D32F71E9D0A368B95795B66F7546F41CA2F0F1C42096D)
, .INIT_27 (256'hAD3A96E180366946521C3AC623510BC8A2188D1777D462584CAE36DF20F70AFF)
, .INIT_28 (256'hC335AA4490DD77115CF2429228040D5AB844A09B888E702E57883EAC25AA0C91)
, .INIT_29 (256'hD8C6BD62A15984C467BC4A592CB60EECCE0CB3DC99217DEE625846762A5D0E23)
, .INIT_2A (256'hEDE2D033B1A7925E727A521C3167107EE364C6D5A9868B956D1D4E3B2F0F0FB5)
, .INIT_2B (256'h027DE2AFC1C19FDC7D2B59DA3617120FF840D97CB9BB992177D455FC33BF1146)
, .INIT_2C (256'h168CF4CFD1A2AD3A87CC61933AC613A10C96EBCBC9B9A68F827D5DB7386F12D8)
, .INIT_2D (256'h2A03068BE146BA76925E69463F741533205BFDBAD97CB3DC8D17656D3D1D146A)
, .INIT_2E (256'h3CDA17DDF0A9C78E9CDF70F2442016C533830F42E900C10797A16D1D41CA15FC)
, .INIT_2F (256'h4F0428BCFFC5D47FA74D789848CB18574605205BF840CE0CA21874C64676178E)
, .INIT_30 (256'h607939230E97E146B1A780364D7519E857D630FF0738DAE8AC7C7C684B20191F)
, .INIT_31 (256'h712F490A1D1AEDE2BBEC87CC521C1B7A68EC412715E3E79AB6CC84024FC91AB1)
, .INIT_32 (256'h811D586B2B4AFA4FC61B8F5B56C21D0B793F50CB243DF41FC1078B95546F1C42)
, .INIT_33 (256'h903A67403923068BD03396E15B661E9D88C65FE732420074CB2A931F59141DD4)
, .INIT_34 (256'h9E7E758246A01294DA329E5D6008202E97776E743FED0C96D5369AA05DB71F65)
, .INIT_35 (256'hABE1832D53BE1E68E418A5D164A821BFA54C7C6B4D3B1885DF28A218625820F7)
, .INIT_36 (256'hB85C903A60792A03EDE2AD3A69462351B23C89C75A28243DE900A98666F72288)
, .INIT_37 (256'hC3E99CA36CCD3565F790B4986DE124E2BE41968366B02FBCF2BDB0EA6B942419)
, .INIT_38 (256'hCE81A86578B7408A0121BBEC727A2673C954A29A72D03AFFFC5DB844702E25AA)
, .INIT_39 (256'hD81EB37A84334B700A94C33577112804D36FAE067E83460505DFBF9274C6273B)
, .INIT_3A (256'hE0BBBDDE8F3E561613E8CA727BA52994DC8DB8C389C750CB0F42C6D5795B28CC)
, .INIT_3B (256'hE853C78C99D560791D1AD1A280362B25E4A8C2CC94985B501885CE0C7DEE2A5D)
, .INIT_3C (256'hEEE3D081A3F46A97262BD8C684C42CB6EBBDCC1E9EF3659121A7D536827D2BEE)
, .INIT_3D (256'hF467D8B9AD98746F2F1ADFDD89502E46F1C7D4B5A8D66F8C2AA7DC53870B2D7E)
, .INIT_3E (256'hF8DBE030B6C07DFD37E4E6E78DD92FD7F6C3DC8DB23C793F3383E3648B952F0F)
, .INIT_3F (256'hFC3EE6E3BF678742408AEDE2925E3167FAAFE3A2BB2482A93C3CEA66901C309F)
, .INITP_00 (256'h5555555555555555555555555555555555555555555555555555555555550001)
, .INITP_01 (256'h5555555555555555555555555555555555555555555555555555555555555555)
, .INITP_02 (256'h1555155555555555555555555555555555555555555555555555555555555555)
, .INITP_03 (256'h0155055505550555055505550555055505550555055515551555155515551555)
, .INITP_04 (256'h0000000000000000000000000000000000000000000000000000000000005540)
, .INITP_05 (256'h5000500050005000500040004000400040000000000000000000000000000000)
, .INITP_06 (256'h5500550055005500550055005500550055005500540054005400540054005400)
, .INITP_07 (256'h5540554055405540554055405540554055405540554055405540554055405500)
