// Created with ./create_bayer_fold_rom.py
// MCLT 16x16...22x22 Bayer -> 8x8 fold indices
, .INIT_00 (256'hA4A4A2A2A6A6A0A0A8A8AEAEAAAAACACB3B3B5B5B1B1B7B7BFBFB9B9BDBDBBBB)
, .INIT_01 (256'h848482828686808088888E8E8A8A8C8C93939595919197979F9F99999D9D9B9B)
, .INIT_02 (256'h13131515111117171F1F19191D1D1B1B040402020606000008080E0E0A0A0C0C)
, .INIT_03 (256'h33333535313137373F3F39393D3D3B3B242422222626202028282E2E2A2A2C2C)
, .INIT_04 (256'hD3D3D5D5D1D1D7D7DFDFD9D9DDDDDBDBC4C4C2C2C6C6C0C0C8C8CECECACACCCC)
, .INIT_05 (256'hF3F3F5F5F1F1F7F7FFFFF9F9FDFDFBFBE4E4E2E2E6E6E0E0E8E8EEEEEAEAECEC)
, .INIT_06 (256'h646462626666606068686E6E6A6A6C6C73737575717177777F7F79797D7D7B7B)
, .INIT_07 (256'h444442424646404048484E4E4A4A4C4C53535555515157575F5F59595D5D5B5B)
, .INIT_08 (256'hA3A3A5A5A1A1A7A7AFAFA9A9ADADABABB4B4B2B2B6B6B0B0B8B8BEBEBABABCBC)
, .INIT_09 (256'h83838585818187878F8F89898D8D8B8B949492929696909098989E9E9A9A9C9C)
, .INIT_0A (256'h141412121616101018181E1E1A1A1C1C03030505010107070F0F09090D0D0B0B)
, .INIT_0B (256'h343432323636303038383E3E3A3A3C3C23232525212127272F2F29292D2D2B2B)
, .INIT_0C (256'hD4D4D2D2D6D6D0D0D8D8DEDEDADADCDCC3C3C5C5C1C1C7C7CFCFC9C9CDCDCBCB)
, .INIT_0D (256'hF4F4F2F2F6F6F0F0F8F8FEFEFAFAFCFCE3E3E5E5E1E1E7E7EFEFE9E9EDEDEBEB)
, .INIT_0E (256'h63636565616167676F6F69696D6D6B6B747472727676707078787E7E7A7A7C7C)
, .INIT_0F (256'h43434545414147474F4F49494D4D4B4B545452525656505058585E5E5A5A5C5C)
, .INIT_10 (256'hB8A4B6A2BAA6B4A0BCA8C2AEBEAAC0ACC9B3CBB5C7B1CDB7D5BFCFB9D3BDD1BB)
, .INIT_11 (256'h948492829686908098889E8E9A8A9C8CA593A795A391A997B19FAB99AF9DAD9B)
, .INIT_12 (256'h1513171513111917211F1B191F1D1D1B040402020606000008080E0E0A0A0C0C)
, .INIT_13 (256'h39333B3537313D37453F3F39433D413B282426222A2624202C28322E2E2A302C)
, .INIT_14 (256'hEDD3EFD5EBD1F1D7F9DFF3D9F7DDF5DBDCC4DAC2DEC6D8C0E0C8E6CEE2CAE4CC)
, .INIT_15 (256'h11F313F50FF115F71DFF17F91BFD19FB00E4FEE202E6FCE004E80AEE06EA08EC)
, .INIT_16 (256'h70646E6272666C6074687A6E766A786C817383757F7185778D7F87798B7D897B)
, .INIT_17 (256'h4C444A424E4648405048564E524A544C5D535F555B516157695F6359675D655B)
, .INIT_18 (256'hB7A3B9A5B5A1BBA7C3AFBDA9C1ADBFABCAB4C8B2CCB6C6B0CEB8D4BED0BAD2BC)
, .INIT_19 (256'h93839585918197879F8F99899D8D9B8BA694A492A896A290AA98B09EAC9AAE9C)
, .INIT_1A (256'h16141412181612101A18201E1C1A1E1C03030505010107070F0F09090D0D0B0B)
, .INIT_1B (256'h3A3438323C3636303E38443E403A423C2723292525212B27332F2D29312D2F2B)
, .INIT_1C (256'hEED4ECD2F0D6EAD0F2D8F8DEF4DAF6DCDBC3DDC5D9C1DFC7E7CFE1C9E5CDE3CB)
, .INIT_1D (256'h12F410F214F60EF016F81CFE18FA1AFCFFE301E5FDE103E70BEF05E909ED07EB)
, .INIT_1E (256'h6F6371656D6173677B6F7569796D776B8274807284767E7086788C7E887A8A7C)
, .INIT_1F (256'h4B434D4549414F47574F5149554D534B5E545C5260565A506258685E645A665C)
, .INIT_20 (256'hCCA4CAA2CEA6C8A0D0A8D6AED2AAD4ACDFB3E1B5DDB1E3B7EBBFE5B9E9BDE7BB)
, .INIT_21 (256'hA484A282A686A080A888AE8EAA8AAC8CB793B995B591BB97C39FBD99C19DBF9B)
, .INIT_22 (256'h1713191515111B17231F1D19211D1F1B040402020606000008080E0E0A0A0C0C)
, .INIT_23 (256'h3F3341353D3143374B3F4539493D473B2C242A222E2628203028362E322A342C)
, .INIT_24 (256'h07D309D505D10BD713DF0DD911DD0FDBF4C4F2C2F6C6F0C0F8C8FECEFACAFCCC)
, .INIT_25 (256'h2FF331F52DF133F73BFF35F939FD37FB1CE41AE21EE618E020E826EE22EA24EC)
, .INIT_26 (256'h7C647A627E6678608068866E826A846C8F7391758D7193779B7F9579997D977B)
, .INIT_27 (256'h544452425646504058485E4E5A4A5C4C6753695565516B57735F6D59715D6F5B)
, .INIT_28 (256'hCBA3CDA5C9A1CFA7D7AFD1A9D5ADD3ABE0B4DEB2E2B6DCB0E4B8EABEE6BAE8BC)
, .INIT_29 (256'hA383A585A181A787AF8FA989AD8DAB8BB894B692BA96B490BC98C29EBE9AC09C)
, .INIT_2A (256'h181416121A1614101C18221E1E1A201C03030505010107070F0F09090D0D0B0B)
, .INIT_2B (256'h40343E3242363C3044384A3E463A483C2B232D2529212F27372F3129352D332B)
, .INIT_2C (256'h08D406D20AD604D00CD812DE0EDA10DCF3C3F5C5F1C1F7C7FFCFF9C9FDCDFBCB)
, .INIT_2D (256'h30F42EF232F62CF034F83AFE36FA38FC1BE31DE519E11FE727EF21E925ED23EB)
, .INIT_2E (256'h7B637D6579617F67876F8169856D836B90748E7292768C7094789A7E967A987C)
, .INIT_2F (256'h53435545514157475F4F59495D4D5B4B685466526A5664506C58725E6E5A705C)
, .INIT_30 (256'hE0A4DEA2E2A6DCA0E4A8EAAEE6AAE8ACF5B3F7B5F3B1F9B701BFFBB9FFBDFDBB)
, .INIT_31 (256'hB484B282B686B080B888BE8EBA8ABC8CC993CB95C791CD97D59FCF99D39DD19B)
, .INIT_32 (256'h19131B1517111D17251F1F19231D211B040402020606000008080E0E0A0A0C0C)
, .INIT_33 (256'h4533473543314937513F4B394F3D4D3B30242E2232262C2034283A2E362A382C)
, .INIT_34 (256'h21D323D51FD125D72DDF27D92BDD29DB0CC40AC20EC608C010C816CE12CA14CC)
, .INIT_35 (256'h4DF34FF54BF151F759FF53F957FD55FB38E436E23AE634E03CE842EE3EEA40EC)
, .INIT_36 (256'h886486628A6684608C68926E8E6A906C9D739F759B71A177A97FA379A77DA57B)
, .INIT_37 (256'h5C445A425E4658406048664E624A644C715373556F5175577D5F77597B5D795B)
, .INIT_38 (256'hDFA3E1A5DDA1E3A7EBAFE5A9E9ADE7ABF6B4F4B2F8B6F2B0FAB800BEFCBAFEBC)
, .INIT_39 (256'hB383B585B181B787BF8FB989BD8DBB8BCA94C892CC96C690CE98D49ED09AD29C)
, .INIT_3A (256'h1A1418121C1616101E18241E201A221C03030505010107070F0F09090D0D0B0B)
, .INIT_3B (256'h46344432483642304A38503E4C3A4E3C2F2331252D2133273B2F3529392D372B)
, .INIT_3C (256'h22D420D224D61ED026D82CDE28DA2ADC0BC30DC509C10FC717CF11C915CD13CB)
, .INIT_3D (256'h4EF44CF250F64AF052F858FE54FA56FC37E339E535E13BE743EF3DE941ED3FEB)
, .INIT_3E (256'h8763896585618B67936F8D69916D8F6B9E749C72A0769A70A278A87EA47AA67C)
, .INIT_3F (256'h5B435D4559415F47674F6149654D634B7254705274566E5076587C5E785A7A5C)
, .INITP_00 (256'hBB88EE22BB88EE22EE22BB88EE22BB8811DD447711DD4477BB88EE22BB88EE22)
, .INITP_01 (256'hEE22BB88EE22BB88BB88EE22BB88EE22447711DD447711DDEE22BB88EE22BB88)
, .INITP_02 (256'hBB88EE22BB88EE22EE22BB88EE22BB8811DD447711DD4477BB88EE22BB88EE22)
, .INITP_03 (256'hEE22BB88EE22BB88BB88EE22BB88EE22447711DD447711DDEE22BB88EE22BB88)
, .INITP_04 (256'hBB88EE22BB88EE22EE22BB88EE22BB8811DD447711DD4477BB88EE22BB88EE22)
, .INITP_05 (256'hEE22BB88EE22BB88BB88EE22BB88EE22447711DD447711DDEE22BB88EE22BB88)
, .INITP_06 (256'hBB88EE22BB88EE22EE22BB88EE22BB8811DD447711DD4477BB88EE22BB88EE22)
, .INITP_07 (256'hEE22BB88EE22BB88BB88EE22BB88EE22447711DD447711DDEE22BB88EE22BB88)
