    parameter FPGA_VERSION =          32'h03930038;