, .INIT_00 (256'h00100000000E0000000C02020035000000220000000C0000000A0000000C0000)
, .INIT_01 (256'h1C3C9449543244190060001B0108001B00500402040401040022000600120000)
, .INIT_02 (256'h001BC8300014000C0210002B2507250E0180001B0003004200180000001B4455)
, .INIT_03 (256'h4C6B2C45141B0012003C01080028000A040800220410001B01020110001B0005)
, .INIT_04 (256'h0210001B14490102005004020404003CB080707D00A0003C8C6E845584C7443A)
, .INIT_05 (256'h000000512507250E0240004F2507250E0240005F0000003C0000001B0210003C)
, .INIT_06 (256'h02200204006E0402009000EEA89968FC18F518D498B058E0388564570C27045B)
, .INIT_07 (256'h003CB0800000005300840022003CB080707D307A30FC02080074D10E5104903C)
, .INIT_08 (256'h2891290A0000000000000014021000892507250E018000A2D1070120003C0000)
, .INIT_09 (256'h0CB6290A0210009D2507250E04400053000C009700050097C895002200440097)
, .INIT_0A (256'h00530081005348AE00220044003C48AE28AA290A0000000000000024003C4882)
, .INIT_0B (256'h0044008800BED1075104042000BA883C08A2003000B6021000B42507250E0240)
, .INIT_0C (256'h0048021000CEC50E2507250700C000C90030003C88A200300009003C88A250C3)
, .INIT_0D (256'h003C34DB000000DD001100DDC8DB021000D82507250E0140003C88A250C30044)
, .INIT_0E (256'h250E0480005301010053C8EC290A0000000000000014021000E42507250E0280)
, .INIT_0F (256'h01002507250E024001020082021000F92507250E0240003C0401021000F22507)
, .INIT_10 (256'h00410410010C0000010C0201010C00210410010C002100840102000001020210)
, .INIT_11 (256'h000000000000000000000000000000000000000000000000000000000000003C)
, .INITP_00 (256'h08802605C240900789C9C8888A000C25062040820809C8020188800222222222)
, .INITP_01 (256'h27209C82720A00270882271A009C86068072E22721816802A89C882068009C32)
, .INITP_02 (256'h0000000000000000000000000000000000000000000000000000000082220822)
