, .INIT_00 (256'h000800F8000700780005001A0004000B0003000400020001000200000004000A)
, .INIT_01 (256'h00020000000000000000000000000000000000000010FF830010FF82000A03F6)
, .INIT_02 (256'h0010FF850010FF84000B07F6000901F6000700790005001B0004000C00000000)
, .INIT_03 (256'h00030002000000000000000000000000000000000010FF880010FF870010FF86)
, .INIT_04 (256'h0010FF8B0010FF8A0010FF89000C0FF4000A03F7000800F90005001C00000000)
, .INIT_05 (256'h00030003000000000000000000000000000000000010FF8E0010FF8D0010FF8C)
, .INIT_06 (256'h0010FF920010FF910010FF900010FF8F000C0FF5000901F70006003A00000000)
, .INIT_07 (256'h00030004000000000000000000000000000000000010FF950010FF940010FF93)
, .INIT_08 (256'h0010FF9A0010FF990010FF980010FF970010FF96000A03F80006003B00000000)
, .INIT_09 (256'h00030005000000000000000000000000000000000010FF9D0010FF9C0010FF9B)
, .INIT_0A (256'h0010FFA20010FFA10010FFA00010FF9F0010FF9E000B07F70007007A00000000)
, .INIT_0B (256'h00030006000000000000000000000000000000000010FFA50010FFA40010FFA3)
, .INIT_0C (256'h0010FFAA0010FFA90010FFA80010FFA70010FFA6000C0FF60007007B00000000)
, .INIT_0D (256'h0004000E000000000000000000000000000000000010FFAD0010FFAC0010FFAB)
, .INIT_0E (256'h0010FFB20010FFB10010FFB00010FFAF0010FFAE000C0FF7000800FA00000000)
, .INIT_0F (256'h0005001E000000000000000000000000000000000010FFB50010FFB40010FFB3)
, .INIT_10 (256'h0010FFBA0010FFB90010FFB80010FFB70010FFB6000F7FC0000901F800000000)
, .INIT_11 (256'h0006003E000000000000000000000000000000000010FFBD0010FFBC0010FFBB)
, .INIT_12 (256'h0010FFC30010FFC20010FFC10010FFC00010FFBF0010FFBE000901F900000000)
, .INIT_13 (256'h0007007E000000000000000000000000000000000010FFC60010FFC50010FFC4)
, .INIT_14 (256'h0010FFCC0010FFCB0010FFCA0010FFC90010FFC80010FFC7000901FA00000000)
, .INIT_15 (256'h000800FE000000000000000000000000000000000010FFCF0010FFCE0010FFCD)
, .INIT_16 (256'h0010FFD50010FFD40010FFD30010FFD20010FFD10010FFD0000A03F900000000)
, .INIT_17 (256'h000901FE000000000000000000000000000000000010FFD80010FFD70010FFD6)
, .INIT_18 (256'h0010FFDE0010FFDD0010FFDC0010FFDB0010FFDA0010FFD9000A03FA00000000)
, .INIT_19 (256'h00000000000000000000000000000000000000000010FFE10010FFE00010FFDF)
, .INIT_1A (256'h0010FFE70010FFE60010FFE50010FFE40010FFE30010FFE2000B07F800000000)
, .INIT_1B (256'h00000000000000000000000000000000000000000010FFEA0010FFE90010FFE8)
, .INIT_1C (256'h0010FFF10010FFF00010FFEF0010FFEE0010FFED0010FFEC0010FFEB00000000)
, .INIT_1D (256'h00000000000000000000000000000000000000000010FFF40010FFF30010FFF2)
, .INIT_1E (256'h0010FFFB0010FFFA0010FFF90010FFF80010FFF70010FFF60010FFF5000B07F9)
, .INIT_1F (256'h00000000000000000000000000000000000000000010FFFE0010FFFD0010FFFC)
, .INIT_20 (256'h000700780006003800050019000500180004000A000300040002000100020000)
, .INIT_21 (256'h0002000000000000000000000000000000000000000C0FF4000A03F6000901F4)
, .INIT_22 (256'h0010FF88000C0FF5000B07F6000901F5000800F6000600390004000B00000000)
, .INIT_23 (256'h00020001000000000000000000000000000000000010FF8B0010FF8A0010FF89)
, .INIT_24 (256'h0010FF8D0010FF8C000F7FC2000C0FF6000A03F7000800F70005001A00000000)
, .INIT_25 (256'h00020002000000000000000000000000000000000010FF900010FF8F0010FF8E)
, .INIT_26 (256'h0010FF930010FF920010FF91000C0FF7000A03F8000800F80005001B00000000)
, .INIT_27 (256'h00030006000000000000000000000000000000000010FF960010FF950010FF94)
, .INIT_28 (256'h0010FF9B0010FF9A0010FF990010FF980010FF97000901F60006003A00000000)
, .INIT_29 (256'h0004000E000000000000000000000000000000000010FF9E0010FF9D0010FF9C)
, .INIT_2A (256'h0010FFA30010FFA20010FFA10010FFA00010FF9F000A03F90006003B00000000)
, .INIT_2B (256'h0005001E000000000000000000000000000000000010FFA60010FFA50010FFA4)
, .INIT_2C (256'h0010FFAB0010FFAA0010FFA90010FFA80010FFA7000B07F70007007900000000)
, .INIT_2D (256'h0006003E000000000000000000000000000000000010FFAE0010FFAD0010FFAC)
, .INIT_2E (256'h0010FFB30010FFB20010FFB10010FFB00010FFAF000B07F80007007A00000000)
, .INIT_2F (256'h0007007E000000000000000000000000000000000010FFB60010FFB50010FFB4)
, .INIT_30 (256'h0010FFBC0010FFBB0010FFBA0010FFB90010FFB80010FFB7000800F900000000)
, .INIT_31 (256'h000800FE000000000000000000000000000000000010FFBF0010FFBE0010FFBD)
, .INIT_32 (256'h0010FFC50010FFC40010FFC30010FFC20010FFC10010FFC0000901F700000000)
, .INIT_33 (256'h000901FE000000000000000000000000000000000010FFC80010FFC70010FFC6)
, .INIT_34 (256'h0010FFCE0010FFCD0010FFCC0010FFCB0010FFCA0010FFC9000901F800000000)
, .INIT_35 (256'h000A03FE000000000000000000000000000000000010FFD10010FFD00010FFCF)
, .INIT_36 (256'h0010FFD70010FFD60010FFD50010FFD40010FFD30010FFD2000901F900000000)
, .INIT_37 (256'h000B07FE000000000000000000000000000000000010FFDA0010FFD90010FFD8)
, .INIT_38 (256'h0010FFE00010FFDF0010FFDE0010FFDD0010FFDC0010FFDB000901FA00000000)
, .INIT_39 (256'h00000000000000000000000000000000000000000010FFE30010FFE20010FFE1)
, .INIT_3A (256'h0010FFE90010FFE80010FFE70010FFE60010FFE50010FFE4000B07F900000000)
, .INIT_3B (256'h00000000000000000000000000000000000000000010FFEC0010FFEB0010FFEA)
, .INIT_3C (256'h0010FFF20010FFF10010FFF00010FFEF0010FFEE0010FFED000E3FE000000000)
, .INIT_3D (256'h00000000000000000000000000000000000000000010FFF50010FFF40010FFF3)
, .INIT_3E (256'h0010FFFB0010FFFA0010FFF90010FFF80010FFF70010FFF6000F7FC3000A03FA)
, .INIT_3F (256'h00000000000000000000000000000000000000000010FFFE0010FFFD0010FFFC)
