, .INIT_00 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_01 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_02 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_03 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_04 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_05 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_06 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_07 (256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
, .INIT_08 (256'h174615551555333340005555800080001555199A200033335555800080005555)
, .INIT_09 (256'h155510000F0F199A2AAB40005555555517461249174620003333555555555555)
, .INIT_0A (256'h0E390B210C31100013B117462492333311110C310BA312491746249240004000)
, .INIT_0B (256'h0CCD0C310CCD0BA30CCD0D790E3912490CCD0AAB0AAB0C310F0F100013B1199A)
, .INIT_0C (256'h0CCD0CCD0CCD0CCD13B13333400040000CCD0CCD0CCD0CCD1C72333340005555)
, .INIT_0D (256'h0CCD0CCD0CCD0CCD0CCD0CCD13B11C720CCD0CCD0CCD0CCD0CCD174633333333)
, .INIT_0E (256'h0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD)
, .INIT_0F (256'h0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD0CCD)
