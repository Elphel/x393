, .INIT_00 (256'h4444444433333333333333332222222222222222111111111111111100000000)
, .INIT_01 (256'h8888888877777777777777776666666666666666555555555555555544444444)
, .INIT_02 (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_03 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_04 (256'h4444444433333333333333332222222222222222111111111111111100000000)
, .INIT_05 (256'h8888888877777777777777776666666666666666555555555555555544444444)
, .INIT_06 (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_07 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_08 (256'h4444444433333333333333322222222222222221111111111111100000000000)
, .INIT_09 (256'h8888888877777777777777776666666666666666555555555555555544444444)
, .INIT_0A (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_0B (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_0C (256'h4444444433333333333333322222222222222221111111111111100000000000)
, .INIT_0D (256'h8888888877777777777777776666666666666666555555555555555544444444)
, .INIT_0E (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_0F (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_10 (256'h4444444333333333333333322222222222222211111111111000000000000000)
, .INIT_11 (256'h8888888877777777777777776666666666666666555555555555555444444444)
, .INIT_12 (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_13 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_14 (256'h4444444333333333333333322222222222222211111111111000000000000000)
, .INIT_15 (256'h8888888877777777777777776666666666666666555555555555555444444444)
, .INIT_16 (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_17 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_18 (256'h4444443333333333333222222222211111111111100000000000000000000000)
, .INIT_19 (256'h8888888877777777777777766666666666666665555555555555555444444444)
, .INIT_1A (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_1B (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_1C (256'h4444443333333333333222222222211111111111100000000000000000000000)
, .INIT_1D (256'h8888888877777777777777766666666666666665555555555555555444444444)
, .INIT_1E (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999988888888)
, .INIT_1F (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_20 (256'h3333333332222222222211111111111111000000000000000000000000000000)
, .INIT_21 (256'h8888888777777777777777766666666666666665555555555555544444444444)
, .INIT_22 (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999888888888)
, .INIT_23 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_24 (256'h3333333332222222222211111111111111000000000000000000000000000000)
, .INIT_25 (256'h8888888777777777777777766666666666666665555555555555544444444444)
, .INIT_26 (256'hCCCCCCCCBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA999999999999999888888888)
, .INIT_27 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_28 (256'h2222222222211111111111111110000000000000000000000000000000000000)
, .INIT_29 (256'h8888888777777777777777666666666666655555555554444444443333333333)
, .INIT_2A (256'hCCCCCCCCBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA9999999999999999888888888)
, .INIT_2B (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_2C (256'h2222222222211111111111111110000000000000000000000000000000000000)
, .INIT_2D (256'h8888888777777777777777666666666666655555555554444444443333333333)
, .INIT_2E (256'hCCCCCCCCBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAA9999999999999999888888888)
, .INIT_2F (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCC)
, .INIT_31 (256'h5555444444443333333333322222222222221111111111111111111111110000)
, .INIT_32 (256'hCCCCCCCBBBBBBBBBBBBBBAAAAAAAAA9999999998888888777777766666665555)
, .INIT_33 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCCC)
, .INIT_35 (256'h5555444444443333333333322222222222221111111111111111111111110000)
, .INIT_36 (256'hCCCCCCCBBBBBBBBBBBBBBAAAAAAAAA9999999998888888777777766666665555)
, .INIT_37 (256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDCCCCCCCCC)
, .INIT_3B (256'hFFFFFFFFFEEDCBA9987766555444333332222222211111111111111111111100)
, .INIT_3F (256'hFFFFFFFFFEEDCBA9987766555444333332222222211111111111111111111100)
