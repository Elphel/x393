, .INITP_00 (INITP_00)
, .INITP_01 (INITP_01)
, .INITP_02 (INITP_02)
, .INITP_03 (INITP_03)
, .INITP_04 (INITP_04)
, .INITP_05 (INITP_05)
, .INITP_06 (INITP_06)
, .INITP_07 (INITP_07)
, .INIT_00  (INIT_00)
, .INIT_01  (INIT_01)
, .INIT_02  (INIT_02)
, .INIT_03  (INIT_03)
, .INIT_04  (INIT_04)
, .INIT_05  (INIT_05)
, .INIT_06  (INIT_06)
, .INIT_07  (INIT_07)
, .INIT_08  (INIT_08)
, .INIT_09  (INIT_09)
, .INIT_0A  (INIT_0A)
, .INIT_0B  (INIT_0B)
, .INIT_0C  (INIT_0C)
, .INIT_0D  (INIT_0D)
, .INIT_0E  (INIT_0E)
, .INIT_0F  (INIT_0F)
, .INIT_10  (INIT_10)
, .INIT_11  (INIT_11)
, .INIT_12  (INIT_12)
, .INIT_13  (INIT_13)
, .INIT_14  (INIT_14)
, .INIT_15  (INIT_15)
, .INIT_16  (INIT_16)
, .INIT_17  (INIT_17)
, .INIT_18  (INIT_18)
, .INIT_19  (INIT_19)
, .INIT_1A  (INIT_1A)
, .INIT_1B  (INIT_1B)
, .INIT_1C  (INIT_1C)
, .INIT_1D  (INIT_1D)
, .INIT_1E  (INIT_1E)
, .INIT_1F  (INIT_1F)
, .INIT_20  (INIT_20)
, .INIT_21  (INIT_21)
, .INIT_22  (INIT_22)
, .INIT_23  (INIT_23)
, .INIT_24  (INIT_24)
, .INIT_25  (INIT_25)
, .INIT_26  (INIT_26)
, .INIT_27  (INIT_27)
, .INIT_28  (INIT_28)
, .INIT_29  (INIT_29)
, .INIT_2A  (INIT_2A)
, .INIT_2B  (INIT_2B)
, .INIT_2C  (INIT_2C)
, .INIT_2D  (INIT_2D)
, .INIT_2E  (INIT_2E)
, .INIT_2F  (INIT_2F)
, .INIT_30  (INIT_30)
, .INIT_31  (INIT_31)
, .INIT_32  (INIT_32)
, .INIT_33  (INIT_33)
, .INIT_34  (INIT_34)
, .INIT_35  (INIT_35)
, .INIT_36  (INIT_36)
, .INIT_37  (INIT_37)
, .INIT_38  (INIT_38)
, .INIT_39  (INIT_39)
, .INIT_3A  (INIT_3A)
, .INIT_3B  (INIT_3B)
, .INIT_3C  (INIT_3C)
, .INIT_3D  (INIT_3D)
, .INIT_3E  (INIT_3E)
, .INIT_3F  (INIT_3F)
